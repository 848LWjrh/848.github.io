module hello_world;
initial begin
	$display("hello_world\n");
end

endmodule
